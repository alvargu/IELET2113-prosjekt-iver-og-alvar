-- Need to fil inn