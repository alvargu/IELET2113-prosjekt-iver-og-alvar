-- library ieee;